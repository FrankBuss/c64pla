library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.all;

entity c64pla7_testbench is
end entity c64pla7_testbench;

architecture test of c64pla7_testbench is

	type Bytes is array (0 to 65535) of std_logic_vector(7 downto 0);
	signal testVectors: Bytes := (
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", x"bf", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", x"fe", x"7f", x"ff", x"7f", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"bf", x"bf", x"bf", x"bf", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", x"ee", x"ee", x"ff", x"ff", 
		x"ee", x"ee", x"ff", x"ff", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", x"cf", x"cf", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", x"df", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", x"fe", x"f7", x"ff", x"f7", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fd", x"fd", x"fd", x"fd", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", x"fb", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", 
		x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff", x"fe", x"fe", x"ff", x"ff"
	);

	signal fe: std_logic := '0';
	signal a13: std_logic := '0';
	signal a14: std_logic := '0';
	signal a15: std_logic := '0';
	signal va14: std_logic := '0';
	signal charen: std_logic := '0';
	signal hiram: std_logic := '0';
	signal loram: std_logic := '0';
	signal cas: std_logic := '0';
	signal romh: std_logic := '0';
	signal roml: std_logic := '0';
	signal io: std_logic := '0';
	signal ramrw: std_logic := '0';
	signal grw: std_logic := '0';
	signal charom: std_logic := '0';
	signal kernal: std_logic := '0';
	signal basic: std_logic := '0';
	signal casram: std_logic := '0';
	signal xoe: std_logic := '0';
	signal va12: std_logic := '0';
	signal va13: std_logic := '0';
	signal game: std_logic := '0';
	signal exrom: std_logic := '0';
	signal rw: std_logic := '0';
	signal aec: std_logic := '0';
	signal ba: std_logic := '0';
	signal a12: std_logic := '0';

begin
	
	c64pla7_inst: entity c64pla7 
		port map(
			fe => fe,
			a13 => a13,
			a14 => a14,
			a15 => a15,
			va14 => va14,
			charen => charen,
			hiram => hiram,
			loram => loram,
			cas => cas,
			romh => romh,
			roml => roml,
			io => io,
			ramrw => ramrw,
			grw => grw,
			charom => charom,
			kernal => kernal,
			basic => basic,
			casram => casram,
			xoe => xoe,
			va12 => va12,
			va13 => va13,
			game => game,
			exrom => exrom,
			rw => rw,
			aec => aec,
			ba => ba,
			a12 => a12
		);

	process
		variable input: std_logic_vector(15 downto 0);
		variable expectedOutput: std_logic_vector(7 downto 0);
		variable i2: integer;
	begin
		xoe <= '0';
		for i in 0 to testVectors'high loop
			i2 := i;
			input := std_logic_vector(to_unsigned(i, input'length));
			cas <= input(1);
			loram <= input(2);
			hiram <= input(3);
			charen <= input(4);
			va14 <= input(5);
			a15 <= input(6);
			a14 <= input(7);
			a13 <= input(12);
			a12 <= input(14);
			ba <= input(13);
			aec <= input(8);
			rw <= input(9);
			exrom <= input(11);
			game <= input(15);
			va13 <= input(10);
			va12 <= input(0);
			wait for 1 ns;
			expectedOutput := testVectors(i);
			assert casram <= expectedOutput(0) report "error" severity failure;
			assert basic <= expectedOutput(1) report "error" severity failure;
			assert kernal <= expectedOutput(2) report "error" severity failure;
			assert charom <= expectedOutput(3) report "error" severity failure;
			assert grw <= expectedOutput(4) report "error" severity failure;
			assert io <= expectedOutput(5) report "error" severity failure;
			assert roml <= expectedOutput(6) report "error" severity failure;
			assert romh <= expectedOutput(7) report "error" severity failure;
		end loop;

		-- show simulation end
		assert false report "no failure, simulation successful" severity failure;
		
	end process;
	

end architecture test;
